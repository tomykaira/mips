-- 110000  000 # fmov
-- 110001  001 # fneg
-- 110010  010 # fadd
-- 110011  011 # fsub
-- 110100  100 # fmul
-- 110101  101 # fmuln
-- 110110  110 # fdiv
-- 110111  111 # fsqrt
